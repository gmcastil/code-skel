library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity top is
    generic (
        PLACEHOLDER     : boolean   := true
    );
    port (
        clk     : in    std_logic;
        rst     : in    std_logic
    );

end entity top;

architecture placeholder of top is

begin

end architecture placeholder;
